`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.12.2021 13:19:46
// Design Name: 
// Module Name: DCT_2D_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module DCT_2D_tb;
     reg [15:0]y0,y1,y2,y3,y4,y5,y6,y7;
     reg [15:0]y8,y9,y10,y11,y12,y13,y14,y15;
     reg [15:0]y16,y17,y18,y19,y20,y21,y22,y23;
     reg [15:0]y24,y25,y26,y27,y28,y29,y30,y31;
     reg [15:0]y32,y33,y34,y35,y36,y37,y38,y39;
     reg [15:0]y40,y41,y42,y43,y44,y45,y46,y47;
     reg [15:0]y48,y49,y50,y51,y52,y53,y54,y55;
     reg [15:0]y56,y57,y58,y59,y60,y61,y62,y63;
     //
     wire [15:0]Y0,Y1,Y2,Y3,Y4,Y5,Y6,Y7;
     wire [15:0]Y8,Y9,Y10,Y11,Y12,Y13,Y14,Y15;
     wire [15:0]Y16,Y17,Y18,Y19,Y20,Y21,Y22,Y23;
     wire [15:0]Y24,Y25,Y26,Y27,Y28,Y29,Y30,Y31;
     wire [15:0]Y32,Y33,Y34,Y35,Y36,Y37,Y38,Y39;
     wire [15:0]Y40,Y41,Y42,Y43,Y44,Y45,Y46,Y47;
     wire [15:0]Y48,Y49,Y50,Y51,Y52,Y53,Y54,Y55;
     wire [15:0]Y56,Y57,Y58,Y59,Y60,Y61,Y62,Y63;
    //
    DCT_2D uut (y0,y1,y2,y3,y4,y5,y6,y7,
      y8,y9,y10,y11,y12,y13,y14,y15,
      y16,y17,y18,y19,y20,y21,y22,y23,
      y24,y25,y26,y27,y28,y29,y30,y31,
      y32,y33,y34,y35,y36,y37,y38,y39,
      y40,y41,y42,y43,y44,y45,y46,y47,
      y48,y49,y50,y51,y52,y53,y54,y55,
      y56,y57,y58,y59,y60,y61,y62,y63,
      Y0,Y1,Y2,Y3,Y4,Y5,Y6,Y7,
      Y8,Y9,Y10,Y11,Y12,Y13,Y14,Y15,
      Y16,Y17,Y18,Y19,Y20,Y21,Y22,Y23,
      Y24,Y25,Y26,Y27,Y28,Y29,Y30,Y31,
      Y32,Y33,Y34,Y35,Y36,Y37,Y38,Y39,
      Y40,Y41,Y42,Y43,Y44,Y45,Y46,Y47,
      Y48,Y49,Y50,Y51,Y52,Y53,Y54,Y55,
      Y56,Y57,Y58,Y59,Y60,Y61,Y62,Y63
    );
        //
        initial
        begin
        y0 = {1'b0,11'b00000010000,4'b0000};  //16
        y1 = {1'b0,11'b00000010100,4'b0000};  //20
        y2 = {1'b0,11'b00000001111,4'b0000};  //15
        y3 = {1'b0,11'b00000011110,4'b0000};  //30
        y4 = {1'b0,11'b00000001100,4'b0000};  //12
        y5 = {1'b0,11'b00000001101,4'b0000};  //13
        y6 = {1'b0,11'b00000001100,4'b0000};  //12
        y7 = {1'b0,11'b00000001101,4'b0000};  //13
        
        y8  = {1'b0,11'b00000010000,4'b0000};  //16
        y9  = {1'b0,11'b00000010100,4'b0000};  //20
        y10 = {1'b0,11'b00000001111,4'b0000};  //15
        y11 = {1'b0,11'b00000011110,4'b0000};  //30
        y12 = {1'b0,11'b00000001100,4'b0000};  //12
        y13 = {1'b0,11'b00000001101,4'b0000};  //13
        y14 = {1'b0,11'b00000001100,4'b0000};  //12
        y15 = {1'b0,11'b00000001101,4'b0000};  //13
        
        y16 = {1'b0,11'b00000010000,4'b0000};  //16
        y17 = {1'b0,11'b00000010100,4'b0000};  //20
        y18 = {1'b0,11'b00000001111,4'b0000};  //15
        y19 = {1'b0,11'b00000011110,4'b0000};  //30
        y20 = {1'b0,11'b00000001100,4'b0000};  //12
        y21 = {1'b0,11'b00000001101,4'b0000};  //13
        y22 = {1'b0,11'b00000001100,4'b0000};  //12
        y23 = {1'b0,11'b00000001101,4'b0000};  //13
        
        y24 = {1'b0,11'b00000010000,4'b0000};  //16
        y25 = {1'b0,11'b00000010100,4'b0000};  //20
        y26 = {1'b0,11'b00000001111,4'b0000};  //15
        y27 = {1'b0,11'b00000011110,4'b0000};  //30
        y28 = {1'b0,11'b00000001100,4'b0000};  //12
        y29 = {1'b0,11'b00000001101,4'b0000};  //13
        y30 = {1'b0,11'b00000001100,4'b0000};  //12
        y31 = {1'b0,11'b00000001101,4'b0000};  //13
        
        y32 = {1'b0,11'b00000010000,4'b0000};  //16
        y33 = {1'b0,11'b00000010100,4'b0000};  //20
        y34 = {1'b0,11'b00000001111,4'b0000};  //15
        y35 = {1'b0,11'b00000011110,4'b0000};  //30
        y36 = {1'b0,11'b00000001100,4'b0000};  //12
        y37 = {1'b0,11'b00000001101,4'b0000};  //13
        y38 = {1'b0,11'b00000001100,4'b0000};  //12
        y39 = {1'b0,11'b00000001101,4'b0000};  //13
        
        y40 = {1'b0,11'b00000010000,4'b0000};  //16
        y41 = {1'b0,11'b00000010100,4'b0000};  //20
        y42 = {1'b0,11'b00000001111,4'b0000};  //15
        y43 = {1'b0,11'b00000011110,4'b0000};  //30
        y44 = {1'b0,11'b00000001100,4'b0000};  //12
        y45 = {1'b0,11'b00000001101,4'b0000};  //13
        y46 = {1'b0,11'b00000001100,4'b0000};  //12
        y47 = {1'b0,11'b00000001101,4'b0000};  //13
        
        y48 = {1'b0,11'b00000010000,4'b0000};  //16
        y49 = {1'b0,11'b00000010100,4'b0000};  //20
        y50 = {1'b0,11'b00000001111,4'b0000};  //15
        y51 = {1'b0,11'b00000011110,4'b0000};  //30
        y52 = {1'b0,11'b00000001100,4'b0000};  //12
        y53 = {1'b0,11'b00000001101,4'b0000};  //13
        y54 = {1'b0,11'b00000001100,4'b0000};  //12
        y55 = {1'b0,11'b00000001101,4'b0000};  //13
        
        y56 = {1'b0,11'b00000010000,4'b0000};  //16
        y57 = {1'b0,11'b00000010100,4'b0000};  //20
        y58 = {1'b0,11'b00000001111,4'b0000};  //15
        y59 = {1'b0,11'b00000011110,4'b0000};  //30
        y60 = {1'b0,11'b00000001100,4'b0000};  //12
        y61 = {1'b0,11'b00000001101,4'b0000};  //13
        y62 = {1'b0,11'b00000001100,4'b0000};  //12
        y63 = {1'b0,11'b00000001101,4'b0000};  //13
        #50;
        end
endmodule

